library ieee;
use ieee.std_logic_1164.all;

entity tb_cont_bin is
end tb_cont_bin;

architecture behav of tb_cont_bin is

	--Declaro componente a testear.
	component cont_bin is 
		port (
				start			:in std_logic;
				clk			:in std_logic;
				reset_low	:in std_logic;
				ok				:out std_logic
				);
		end component;
		
	--Señales test bench:
	signal start_tb 		:std_logic := '0';
	signal clk_tb			:std_logic := '0';
	signal reset_low_tb	:std_logic := '0';
	signal ok_tb				:std_logic;
				
	constant clk_semiperiod : time := 50 us;			
				
begin

	uut: cont_bin port map (start => start_tb, clk => clk_tb, reset_low => reset_low_tb, ok => ok_tb);

	clk_tb <= not clk_tb after clk_semiperiod;
	
	data_gen: process 
		begin 
			
			--El reset se encuentra habilitado por lo tanto la salida es un nivel logico bajo.
			wait until clk_tb = '1';
			
			--Desahilitamos el reset y habilitamos start para que comienze a operar el contador.
			reset_low_tb <= '1';
			start_tb <= '1';
			wait until clk_tb = '1';
			
			--Esperamos 11 periodos para observar la salida.
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			wait until clk_tb = '1';
			
			--Luego reseteamos el contador para llevar la salida a cero logico.
			reset_low_tb <= '0';
			wait until clk_tb = '1';
			
		end process;	
			
	
end behav;